
package ahb_apb_pkg;

    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    `include "ahb_xtn.sv"
    `include "apb_xtn.sv"
    `include "ahb_config.sv"
    `include "apb_config.sv"
    `include "ahb_apb_env_config.sv"
    
    `include "ahb_driver.sv"
    `include "ahb_monitor.sv"
    `include "ahb_seqr.sv"
    `include "ahb_agent.sv"
    `include "ahb_top.sv"
    `include "ahb_seq.sv"
    
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_seqr.sv"
    `include "apb_agent.sv"
    `include "apb_top.sv"
    `include "apb_seq.sv"
    
    `include "ahb_apb_virtual_seqr.sv"
    `include "ahb_apb_virtual_seq.sv"
    `include "ahb_apb_scoreboard.sv"
    `include "ahb_apb_env.sv"
    
    `include "ahb_apb_test.sv"

endpackage
